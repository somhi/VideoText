library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"d8d1c187",
    12 => x"48c0c84e",
    13 => x"d5c128c2",
    14 => x"ead6e5ea",
    15 => x"c1467149",
    16 => x"87f90188",
    17 => x"49d8d1c1",
    18 => x"48cccdc1",
    19 => x"0389d089",
    20 => x"404040c0",
    21 => x"d087f640",
    22 => x"50c00581",
    23 => x"f90589c1",
    24 => x"c9cdc187",
    25 => x"c5cdc14d",
    26 => x"02ad744c",
    27 => x"0f2487c4",
    28 => x"c2dc87f7",
    29 => x"c9cdc187",
    30 => x"c9cdc14d",
    31 => x"02ad744c",
    32 => x"8cc487c6",
    33 => x"87f50f6c",
    34 => x"1e87fd00",
    35 => x"4a7186fc",
    36 => x"6949c0ff",
    37 => x"98c0c448",
    38 => x"98487e70",
    39 => x"7287f402",
    40 => x"8efc4879",
    41 => x"731e4f26",
    42 => x"a9738148",
    43 => x"1287c502",
    44 => x"87f60553",
    45 => x"ff1e4f26",
    46 => x"ffc348d4",
    47 => x"26486878",
    48 => x"d4ff1e4f",
    49 => x"78ffc348",
    50 => x"c048d0ff",
    51 => x"d4ff78e1",
    52 => x"2678d448",
    53 => x"d0ff1e4f",
    54 => x"78e0c048",
    55 => x"ff1e4f26",
    56 => x"497087d4",
    57 => x"87c60299",
    58 => x"05a9fbc0",
    59 => x"487187f1",
    60 => x"5e0e4f26",
    61 => x"710e5c5b",
    62 => x"fe4cc04b",
    63 => x"497087f8",
    64 => x"f9c00299",
    65 => x"a9ecc087",
    66 => x"87f2c002",
    67 => x"02a9fbc0",
    68 => x"cc87ebc0",
    69 => x"03acb766",
    70 => x"66d087c7",
    71 => x"7187c202",
    72 => x"02997153",
    73 => x"84c187c2",
    74 => x"7087cbfe",
    75 => x"cd029949",
    76 => x"a9ecc087",
    77 => x"c087c702",
    78 => x"ff05a9fb",
    79 => x"66d087d5",
    80 => x"c087c302",
    81 => x"ecc07b97",
    82 => x"87c405a9",
    83 => x"87c54a74",
    84 => x"0ac04a74",
    85 => x"2648728a",
    86 => x"264b264c",
    87 => x"d5fd1e4f",
    88 => x"4a497087",
    89 => x"04aaf0c0",
    90 => x"f9c087c9",
    91 => x"87c301aa",
    92 => x"c18af0c0",
    93 => x"c904aac1",
    94 => x"aadac187",
    95 => x"c087c301",
    96 => x"48728af7",
    97 => x"261e4f26",
    98 => x"4f261e4f",
    99 => x"1e4f261e",
   100 => x"f8c049c0",
   101 => x"4f2687eb",
   102 => x"494a711e",
   103 => x"dcdf91cc",
   104 => x"c181c881",
   105 => x"1148d0cd",
   106 => x"a2f0c050",
   107 => x"87dbfb49",
   108 => x"ded649c0",
   109 => x"1e4f2687",
   110 => x"c34ad4ff",
   111 => x"d0ff7aff",
   112 => x"78e1c048",
   113 => x"7a717ade",
   114 => x"28b7c848",
   115 => x"48717a70",
   116 => x"7028b7d0",
   117 => x"d848717a",
   118 => x"7a7028b7",
   119 => x"c048d0ff",
   120 => x"4f2678e0",
   121 => x"5c5b5e0e",
   122 => x"86f40e5d",
   123 => x"cc494d71",
   124 => x"81dcdf91",
   125 => x"ca4aa1c8",
   126 => x"a6c47ea1",
   127 => x"cccdc148",
   128 => x"976e78bf",
   129 => x"66c44bbf",
   130 => x"122c734c",
   131 => x"58a6cc48",
   132 => x"84c19c70",
   133 => x"699781c9",
   134 => x"04acb749",
   135 => x"4cc087c2",
   136 => x"4abf976e",
   137 => x"724966c8",
   138 => x"c4b9ff31",
   139 => x"48749966",
   140 => x"4a703072",
   141 => x"d0cdc1b1",
   142 => x"fafd7159",
   143 => x"c11ec787",
   144 => x"1ebfd4cd",
   145 => x"c11edcdf",
   146 => x"bf97d0cd",
   147 => x"87f3c149",
   148 => x"f4c04975",
   149 => x"8ee887ca",
   150 => x"4c264d26",
   151 => x"4f264b26",
   152 => x"711e731e",
   153 => x"fbfd494b",
   154 => x"fd497387",
   155 => x"4b2687f6",
   156 => x"731e4f26",
   157 => x"c24b711e",
   158 => x"d6024aa3",
   159 => x"058ac187",
   160 => x"c187e2c0",
   161 => x"02bfd4cd",
   162 => x"c14887db",
   163 => x"d8cdc188",
   164 => x"c187d258",
   165 => x"02bfd8cd",
   166 => x"cdc187cb",
   167 => x"c148bfd4",
   168 => x"d8cdc180",
   169 => x"c11ec758",
   170 => x"1ebfd4cd",
   171 => x"c11edcdf",
   172 => x"bf97d0cd",
   173 => x"7387cc49",
   174 => x"e3f2c049",
   175 => x"268ef487",
   176 => x"0e4f264b",
   177 => x"5d5c5b5e",
   178 => x"86ccff0e",
   179 => x"59a6e4c0",
   180 => x"c048a6cc",
   181 => x"c080c478",
   182 => x"c180c478",
   183 => x"c47866c8",
   184 => x"c478c180",
   185 => x"c178c180",
   186 => x"c148d8cd",
   187 => x"87d1f778",
   188 => x"f787ebf7",
   189 => x"4c7087c0",
   190 => x"02acfbc0",
   191 => x"c087efc1",
   192 => x"c10566e0",
   193 => x"c4c187e5",
   194 => x"82c44a66",
   195 => x"f4dc7e6a",
   196 => x"20496e48",
   197 => x"10412041",
   198 => x"66c4c151",
   199 => x"78c6c648",
   200 => x"81c7496a",
   201 => x"c4c15174",
   202 => x"81c84966",
   203 => x"a6d851c1",
   204 => x"c178c248",
   205 => x"c94966c4",
   206 => x"c151c081",
   207 => x"ca4966c4",
   208 => x"c151c081",
   209 => x"6a1ed81e",
   210 => x"f681c849",
   211 => x"86c887e4",
   212 => x"4866c8c1",
   213 => x"c701a8c0",
   214 => x"48a6d087",
   215 => x"87ce78c1",
   216 => x"4866c8c1",
   217 => x"a6d888c1",
   218 => x"f587c358",
   219 => x"9c7487f0",
   220 => x"87c0cd02",
   221 => x"c14866d0",
   222 => x"03a866cc",
   223 => x"c887f5cc",
   224 => x"78c048a6",
   225 => x"87eef47e",
   226 => x"d0c14c70",
   227 => x"e2c205ac",
   228 => x"48a6c487",
   229 => x"c4f7786e",
   230 => x"487e7087",
   231 => x"06a866cc",
   232 => x"a6cc87c5",
   233 => x"f4786e48",
   234 => x"4c7087cc",
   235 => x"05acecc0",
   236 => x"d087eac1",
   237 => x"91cc4966",
   238 => x"8166c4c1",
   239 => x"6a4aa1c4",
   240 => x"4aa1c84d",
   241 => x"d8c6526e",
   242 => x"87eaf379",
   243 => x"029c4c70",
   244 => x"fbc087d8",
   245 => x"87d202ac",
   246 => x"d9f35574",
   247 => x"9c4c7087",
   248 => x"c087c702",
   249 => x"ff05acfb",
   250 => x"e0c087ee",
   251 => x"55c1c255",
   252 => x"c07d97c0",
   253 => x"c44866e0",
   254 => x"db05a866",
   255 => x"4866d087",
   256 => x"04a866d4",
   257 => x"66d087ca",
   258 => x"d480c148",
   259 => x"87c858a6",
   260 => x"c14866d4",
   261 => x"58a6d888",
   262 => x"7087dbf2",
   263 => x"acd0c14c",
   264 => x"dc87c905",
   265 => x"80c14866",
   266 => x"58a6e0c0",
   267 => x"02acd0c1",
   268 => x"6e87defd",
   269 => x"66e0c048",
   270 => x"d8c905a8",
   271 => x"a6e4c087",
   272 => x"7478c048",
   273 => x"88fbc048",
   274 => x"7058a6c8",
   275 => x"c9c90298",
   276 => x"88cb4887",
   277 => x"7058a6c8",
   278 => x"ccc10298",
   279 => x"88c94887",
   280 => x"7058a6c8",
   281 => x"f6c30298",
   282 => x"88c44887",
   283 => x"7058a6c8",
   284 => x"87cf0298",
   285 => x"c888c148",
   286 => x"987058a6",
   287 => x"87dfc302",
   288 => x"c887cac8",
   289 => x"f0c048a6",
   290 => x"87eaf078",
   291 => x"ecc04c70",
   292 => x"87c302ac",
   293 => x"c05ca6cc",
   294 => x"cc02acec",
   295 => x"87d6f087",
   296 => x"ecc04c70",
   297 => x"f4ff05ac",
   298 => x"acecc087",
   299 => x"f087c302",
   300 => x"1ec087c4",
   301 => x"66d81eca",
   302 => x"c191cc49",
   303 => x"714866cc",
   304 => x"58a6cc80",
   305 => x"c44866c8",
   306 => x"58a6d080",
   307 => x"49bf66cc",
   308 => x"c187dff0",
   309 => x"d41ede1e",
   310 => x"f049bf66",
   311 => x"86d087d4",
   312 => x"c0484970",
   313 => x"ecc08808",
   314 => x"a8c058a6",
   315 => x"87eec006",
   316 => x"4866e8c0",
   317 => x"c003a8dd",
   318 => x"66c487e4",
   319 => x"e8c049bf",
   320 => x"e0c08166",
   321 => x"66e8c051",
   322 => x"c481c149",
   323 => x"c281bf66",
   324 => x"e8c051c1",
   325 => x"81c24966",
   326 => x"81bf66c4",
   327 => x"486e51c0",
   328 => x"6e78c6c6",
   329 => x"d881c849",
   330 => x"496e5166",
   331 => x"66dc81c9",
   332 => x"ca496e51",
   333 => x"5166c881",
   334 => x"c14866d8",
   335 => x"58a6dc80",
   336 => x"d44866d0",
   337 => x"cb04a866",
   338 => x"4866d087",
   339 => x"a6d480c1",
   340 => x"87c6c558",
   341 => x"c14866d4",
   342 => x"58a6d888",
   343 => x"ef87fbc4",
   344 => x"ecc087fb",
   345 => x"f4ef58a6",
   346 => x"a6f0c087",
   347 => x"a8ecc058",
   348 => x"87c9c005",
   349 => x"e8c048a6",
   350 => x"c3c07866",
   351 => x"87f6ec87",
   352 => x"cc4966d0",
   353 => x"66c4c191",
   354 => x"c8807148",
   355 => x"66c458a6",
   356 => x"c482c84a",
   357 => x"81ca4966",
   358 => x"5166e8c0",
   359 => x"4966ecc0",
   360 => x"e8c081c1",
   361 => x"48c18966",
   362 => x"49703071",
   363 => x"977189c1",
   364 => x"cccdc17a",
   365 => x"e8c049bf",
   366 => x"6a972966",
   367 => x"9871484a",
   368 => x"58a6f4c0",
   369 => x"c44866c4",
   370 => x"58a6cc80",
   371 => x"4dbf66c8",
   372 => x"4866e0c0",
   373 => x"c002a86e",
   374 => x"7ec087c5",
   375 => x"c187c2c0",
   376 => x"c01e6e7e",
   377 => x"49751ee0",
   378 => x"c887c7ec",
   379 => x"c04c7086",
   380 => x"c106acb7",
   381 => x"857487d1",
   382 => x"49bf66c8",
   383 => x"7581e0c0",
   384 => x"c0dd4b89",
   385 => x"ddea714a",
   386 => x"7585c287",
   387 => x"66e4c07e",
   388 => x"c080c148",
   389 => x"c058a6e8",
   390 => x"c14966f0",
   391 => x"02a97081",
   392 => x"c087c5c0",
   393 => x"87c2c04d",
   394 => x"1e754dc1",
   395 => x"49bf66cc",
   396 => x"c481e0c0",
   397 => x"1e718966",
   398 => x"ea4966c8",
   399 => x"86c887f4",
   400 => x"01a8b7c0",
   401 => x"c087c6ff",
   402 => x"c00266e4",
   403 => x"66c487d2",
   404 => x"c081c949",
   405 => x"c45166e4",
   406 => x"e4c74866",
   407 => x"87cdc078",
   408 => x"c94966c4",
   409 => x"c451c281",
   410 => x"e0c94866",
   411 => x"4866d078",
   412 => x"04a866d4",
   413 => x"d087cbc0",
   414 => x"80c14866",
   415 => x"c058a6d4",
   416 => x"66d487d8",
   417 => x"d888c148",
   418 => x"cdc058a6",
   419 => x"87cee987",
   420 => x"c5c04c70",
   421 => x"87c6e987",
   422 => x"66dc4c70",
   423 => x"c080c148",
   424 => x"7458a6e0",
   425 => x"cbc0029c",
   426 => x"4866d087",
   427 => x"a866ccc1",
   428 => x"87cbf304",
   429 => x"c74866d0",
   430 => x"e1c003a8",
   431 => x"4c66d087",
   432 => x"48d8cdc1",
   433 => x"497478c0",
   434 => x"c4c191cc",
   435 => x"a1c48166",
   436 => x"c04a6a4a",
   437 => x"84c17952",
   438 => x"ff04acc7",
   439 => x"e0c087e2",
   440 => x"e0c00266",
   441 => x"66c4c187",
   442 => x"81d4c149",
   443 => x"4a66c4c1",
   444 => x"c082dcc1",
   445 => x"79d8c652",
   446 => x"4966c4c1",
   447 => x"dd81d8c1",
   448 => x"d4c079c4",
   449 => x"66c4c187",
   450 => x"81d4c149",
   451 => x"4a66c4c1",
   452 => x"dd82d8c1",
   453 => x"cfc67acc",
   454 => x"66c4c179",
   455 => x"81e0c149",
   456 => x"e679f2c9",
   457 => x"66cc87ef",
   458 => x"8eccff48",
   459 => x"4c264d26",
   460 => x"4f264b26",
   461 => x"64616f4c",
   462 => x"202e2a20",
   463 => x"00000000",
   464 => x"0000203a",
   465 => x"61422080",
   466 => x"00006b63",
   467 => x"78452080",
   468 => x"1e007469",
   469 => x"cdc11ec7",
   470 => x"df1ebfd4",
   471 => x"cdc11edc",
   472 => x"49bf97d0",
   473 => x"df87dced",
   474 => x"e1c049dc",
   475 => x"8ef487c0",
   476 => x"c01e4f26",
   477 => x"1e4f2648",
   478 => x"c087fac6",
   479 => x"df48f4e0",
   480 => x"e8fe78d0",
   481 => x"e0c049a0",
   482 => x"49c787e4",
   483 => x"c187d1df",
   484 => x"ece0c049",
   485 => x"48d4ff87",
   486 => x"c178ffc3",
   487 => x"c048d4cd",
   488 => x"d0cdc178",
   489 => x"4950c048",
   490 => x"ff87e8fe",
   491 => x"4a7087c4",
   492 => x"87cb029a",
   493 => x"5af8e0c0",
   494 => x"e3de49c7",
   495 => x"c087c587",
   496 => x"87fddf49",
   497 => x"c087e8c2",
   498 => x"fa87dee1",
   499 => x"004f2687",
   500 => x"746f6f42",
   501 => x"2e676e69",
   502 => x"00002e2e",
   503 => x"00000189",
   504 => x"0000135c",
   505 => x"00000000",
   506 => x"00000189",
   507 => x"0000137a",
   508 => x"00000000",
   509 => x"00000189",
   510 => x"00001398",
   511 => x"00000000",
   512 => x"00000189",
   513 => x"000013b6",
   514 => x"00000000",
   515 => x"00000189",
   516 => x"000013d4",
   517 => x"00000000",
   518 => x"00000189",
   519 => x"000013f2",
   520 => x"00000000",
   521 => x"00000189",
   522 => x"00001410",
   523 => x"00000000",
   524 => x"00000198",
   525 => x"00000000",
   526 => x"00000000",
   527 => x"0000018c",
   528 => x"00000000",
   529 => x"00000000",
   530 => x"db86fc1e",
   531 => x"fc7e7087",
   532 => x"1e4f268e",
   533 => x"c048f0fe",
   534 => x"7909cd78",
   535 => x"1e4f2609",
   536 => x"49c8e1c0",
   537 => x"4f2687ed",
   538 => x"bff0fe1e",
   539 => x"1e4f2648",
   540 => x"c148f0fe",
   541 => x"1e4f2678",
   542 => x"c048f0fe",
   543 => x"1e4f2678",
   544 => x"52c04a71",
   545 => x"0e4f2651",
   546 => x"5d5c5b5e",
   547 => x"7186f40e",
   548 => x"7e6d974d",
   549 => x"974ca5c1",
   550 => x"a6c8486c",
   551 => x"c4486e58",
   552 => x"c505a866",
   553 => x"c048ff87",
   554 => x"caff87e6",
   555 => x"49a5c287",
   556 => x"714b6c97",
   557 => x"6b974ba3",
   558 => x"7e6c974b",
   559 => x"80c1486e",
   560 => x"c758a6c8",
   561 => x"58a6cc98",
   562 => x"fe7c9770",
   563 => x"487387e1",
   564 => x"4d268ef4",
   565 => x"4b264c26",
   566 => x"5e0e4f26",
   567 => x"f40e5c5b",
   568 => x"d84c7186",
   569 => x"ffc34a66",
   570 => x"4ba4c29a",
   571 => x"73496c97",
   572 => x"517249a1",
   573 => x"6e7e6c97",
   574 => x"c880c148",
   575 => x"98c758a6",
   576 => x"7058a6cc",
   577 => x"268ef454",
   578 => x"264b264c",
   579 => x"86fc1e4f",
   580 => x"e087e4fd",
   581 => x"c0494abf",
   582 => x"0299c0e0",
   583 => x"1e7287cb",
   584 => x"49f0d0c1",
   585 => x"c487f3fe",
   586 => x"87fcfc86",
   587 => x"fefc7e70",
   588 => x"268efc87",
   589 => x"d0c11e4f",
   590 => x"c2fd49f0",
   591 => x"cde4c087",
   592 => x"87cffc49",
   593 => x"2687edc3",
   594 => x"5b5e0e4f",
   595 => x"fc0e5d5c",
   596 => x"ff7e7186",
   597 => x"d0c14dd4",
   598 => x"eafc49f0",
   599 => x"c04b7087",
   600 => x"c204abb7",
   601 => x"f0c387f8",
   602 => x"87c905ab",
   603 => x"48ece8c0",
   604 => x"d9c278c1",
   605 => x"abe0c387",
   606 => x"c087c905",
   607 => x"c148f0e8",
   608 => x"87cac278",
   609 => x"bff0e8c0",
   610 => x"c287c602",
   611 => x"c24ca3c0",
   612 => x"c04c7387",
   613 => x"02bfece8",
   614 => x"7487e0c0",
   615 => x"29b7c449",
   616 => x"c8eac091",
   617 => x"cf4a7481",
   618 => x"c192c29a",
   619 => x"70307248",
   620 => x"72baff4a",
   621 => x"70986948",
   622 => x"7487db79",
   623 => x"29b7c449",
   624 => x"c8eac091",
   625 => x"cf4a7481",
   626 => x"c392c29a",
   627 => x"70307248",
   628 => x"b069484a",
   629 => x"056e7970",
   630 => x"ff87e7c0",
   631 => x"e1c848d0",
   632 => x"c07dc578",
   633 => x"02bff0e8",
   634 => x"e0c387c3",
   635 => x"ece8c07d",
   636 => x"87c302bf",
   637 => x"737df0c3",
   638 => x"48d0ff7d",
   639 => x"c078e1c8",
   640 => x"e8c078e0",
   641 => x"78c048f0",
   642 => x"48ece8c0",
   643 => x"d0c178c0",
   644 => x"f2f949f0",
   645 => x"c04b7087",
   646 => x"fd03abb7",
   647 => x"48c087c8",
   648 => x"4d268efc",
   649 => x"4b264c26",
   650 => x"00004f26",
   651 => x"00000000",
   652 => x"00000000",
   653 => x"724ac01e",
   654 => x"c091c449",
   655 => x"c081c8ea",
   656 => x"d082c179",
   657 => x"ee04aab7",
   658 => x"0e4f2687",
   659 => x"5d5c5b5e",
   660 => x"f84d710e",
   661 => x"4a7587e1",
   662 => x"922ab7c4",
   663 => x"82c8eac0",
   664 => x"9ccf4c75",
   665 => x"496a94c2",
   666 => x"c32b744b",
   667 => x"7448c29b",
   668 => x"ff4c7030",
   669 => x"714874bc",
   670 => x"f77a7098",
   671 => x"487387f1",
   672 => x"4c264d26",
   673 => x"4f264b26",
   674 => x"00000000",
   675 => x"00000000",
   676 => x"00000000",
   677 => x"00000000",
   678 => x"00000000",
   679 => x"00000000",
   680 => x"00000000",
   681 => x"00000000",
   682 => x"00000000",
   683 => x"00000000",
   684 => x"00000000",
   685 => x"00000000",
   686 => x"00000000",
   687 => x"00000000",
   688 => x"00000000",
   689 => x"00000000",
   690 => x"48d0ff1e",
   691 => x"7178e1c8",
   692 => x"08d4ff48",
   693 => x"4866c478",
   694 => x"7808d4ff",
   695 => x"711e4f26",
   696 => x"4966c44a",
   697 => x"ff49721e",
   698 => x"d0ff87de",
   699 => x"78e0c048",
   700 => x"4f268efc",
   701 => x"711e731e",
   702 => x"4966c84b",
   703 => x"c14a731e",
   704 => x"ff49a2e0",
   705 => x"8efc87d8",
   706 => x"4f264b26",
   707 => x"48d0ff1e",
   708 => x"7178c9c8",
   709 => x"08d4ff48",
   710 => x"1e4f2678",
   711 => x"eb494a71",
   712 => x"48d0ff87",
   713 => x"4f2678c8",
   714 => x"711e731e",
   715 => x"c8d1c14b",
   716 => x"87c302bf",
   717 => x"ff87ebc2",
   718 => x"c9c848d0",
   719 => x"c0487378",
   720 => x"d4ffb0e0",
   721 => x"d0c17808",
   722 => x"78c048fc",
   723 => x"c50266c8",
   724 => x"49ffc387",
   725 => x"49c087c2",
   726 => x"59c4d1c1",
   727 => x"c60266cc",
   728 => x"d5d5c587",
   729 => x"cf87c44a",
   730 => x"c14affff",
   731 => x"c15ac8d1",
   732 => x"c148c8d1",
   733 => x"264b2678",
   734 => x"5b5e0e4f",
   735 => x"710e5d5c",
   736 => x"c4d1c14d",
   737 => x"9d754bbf",
   738 => x"4987cb02",
   739 => x"ecc091c8",
   740 => x"82714ae0",
   741 => x"f0c087c4",
   742 => x"4cc04ae0",
   743 => x"99734912",
   744 => x"bfc0d1c1",
   745 => x"ffb87148",
   746 => x"c17808d4",
   747 => x"c8842bb7",
   748 => x"e704acb7",
   749 => x"fcd0c187",
   750 => x"80c848bf",
   751 => x"58c0d1c1",
   752 => x"4c264d26",
   753 => x"4f264b26",
   754 => x"711e731e",
   755 => x"9a4a134b",
   756 => x"7287cb02",
   757 => x"87e1fe49",
   758 => x"059a4a13",
   759 => x"4b2687f5",
   760 => x"c11e4f26",
   761 => x"49bffcd0",
   762 => x"48fcd0c1",
   763 => x"c478a1c1",
   764 => x"03a9b7c0",
   765 => x"d4ff87db",
   766 => x"c0d1c148",
   767 => x"d0c178bf",
   768 => x"c149bffc",
   769 => x"c148fcd0",
   770 => x"c0c478a1",
   771 => x"e504a9b7",
   772 => x"48d0ff87",
   773 => x"d1c178c8",
   774 => x"78c048c8",
   775 => x"00004f26",
   776 => x"00000000",
   777 => x"00000000",
   778 => x"5f000000",
   779 => x"0000005f",
   780 => x"00030300",
   781 => x"00000303",
   782 => x"147f7f14",
   783 => x"00147f7f",
   784 => x"6b2e2400",
   785 => x"00123a6b",
   786 => x"18366a4c",
   787 => x"0032566c",
   788 => x"594f7e30",
   789 => x"40683a77",
   790 => x"07040000",
   791 => x"00000003",
   792 => x"3e1c0000",
   793 => x"00004163",
   794 => x"63410000",
   795 => x"00001c3e",
   796 => x"1c3e2a08",
   797 => x"082a3e1c",
   798 => x"3e080800",
   799 => x"0008083e",
   800 => x"e0800000",
   801 => x"00000060",
   802 => x"08080800",
   803 => x"00080808",
   804 => x"60000000",
   805 => x"00000060",
   806 => x"18306040",
   807 => x"0103060c",
   808 => x"597f3e00",
   809 => x"003e7f4d",
   810 => x"7f060400",
   811 => x"0000007f",
   812 => x"71634200",
   813 => x"00464f59",
   814 => x"49632200",
   815 => x"00367f49",
   816 => x"13161c18",
   817 => x"00107f7f",
   818 => x"45672700",
   819 => x"00397d45",
   820 => x"4b7e3c00",
   821 => x"00307949",
   822 => x"71010100",
   823 => x"00070f79",
   824 => x"497f3600",
   825 => x"00367f49",
   826 => x"494f0600",
   827 => x"001e3f69",
   828 => x"66000000",
   829 => x"00000066",
   830 => x"e6800000",
   831 => x"00000066",
   832 => x"14080800",
   833 => x"00222214",
   834 => x"14141400",
   835 => x"00141414",
   836 => x"14222200",
   837 => x"00080814",
   838 => x"51030200",
   839 => x"00060f59",
   840 => x"5d417f3e",
   841 => x"001e1f55",
   842 => x"097f7e00",
   843 => x"007e7f09",
   844 => x"497f7f00",
   845 => x"00367f49",
   846 => x"633e1c00",
   847 => x"00414141",
   848 => x"417f7f00",
   849 => x"001c3e63",
   850 => x"497f7f00",
   851 => x"00414149",
   852 => x"097f7f00",
   853 => x"00010109",
   854 => x"417f3e00",
   855 => x"007a7b49",
   856 => x"087f7f00",
   857 => x"007f7f08",
   858 => x"7f410000",
   859 => x"0000417f",
   860 => x"40602000",
   861 => x"003f7f40",
   862 => x"1c087f7f",
   863 => x"00416336",
   864 => x"407f7f00",
   865 => x"00404040",
   866 => x"0c067f7f",
   867 => x"007f7f06",
   868 => x"0c067f7f",
   869 => x"007f7f18",
   870 => x"417f3e00",
   871 => x"003e7f41",
   872 => x"097f7f00",
   873 => x"00060f09",
   874 => x"61417f3e",
   875 => x"00407e7f",
   876 => x"097f7f00",
   877 => x"00667f19",
   878 => x"4d6f2600",
   879 => x"00327b59",
   880 => x"7f010100",
   881 => x"0001017f",
   882 => x"407f3f00",
   883 => x"003f7f40",
   884 => x"703f0f00",
   885 => x"000f3f70",
   886 => x"18307f7f",
   887 => x"007f7f30",
   888 => x"1c366341",
   889 => x"4163361c",
   890 => x"7c060301",
   891 => x"0103067c",
   892 => x"4d597161",
   893 => x"00414347",
   894 => x"7f7f0000",
   895 => x"00004141",
   896 => x"0c060301",
   897 => x"40603018",
   898 => x"41410000",
   899 => x"00007f7f",
   900 => x"03060c08",
   901 => x"00080c06",
   902 => x"80808080",
   903 => x"00808080",
   904 => x"03000000",
   905 => x"00000407",
   906 => x"54742000",
   907 => x"00787c54",
   908 => x"447f7f00",
   909 => x"00387c44",
   910 => x"447c3800",
   911 => x"00004444",
   912 => x"447c3800",
   913 => x"007f7f44",
   914 => x"547c3800",
   915 => x"00185c54",
   916 => x"7f7e0400",
   917 => x"00000505",
   918 => x"a4bc1800",
   919 => x"007cfca4",
   920 => x"047f7f00",
   921 => x"00787c04",
   922 => x"3d000000",
   923 => x"0000407d",
   924 => x"80808000",
   925 => x"00007dfd",
   926 => x"107f7f00",
   927 => x"00446c38",
   928 => x"3f000000",
   929 => x"0000407f",
   930 => x"180c7c7c",
   931 => x"00787c0c",
   932 => x"047c7c00",
   933 => x"00787c04",
   934 => x"447c3800",
   935 => x"00387c44",
   936 => x"24fcfc00",
   937 => x"00183c24",
   938 => x"243c1800",
   939 => x"00fcfc24",
   940 => x"047c7c00",
   941 => x"00080c04",
   942 => x"545c4800",
   943 => x"00207454",
   944 => x"7f3f0400",
   945 => x"00004444",
   946 => x"407c3c00",
   947 => x"007c7c40",
   948 => x"603c1c00",
   949 => x"001c3c60",
   950 => x"30607c3c",
   951 => x"003c7c60",
   952 => x"10386c44",
   953 => x"00446c38",
   954 => x"e0bc1c00",
   955 => x"001c3c60",
   956 => x"74644400",
   957 => x"00444c5c",
   958 => x"3e080800",
   959 => x"00414177",
   960 => x"7f000000",
   961 => x"0000007f",
   962 => x"77414100",
   963 => x"0008083e",
   964 => x"03010102",
   965 => x"00010202",
   966 => x"7f7f7f7f",
   967 => x"007f7f7f",
   968 => x"1c1c0808",
   969 => x"7f7f3e3e",
   970 => x"3e3e7f7f",
   971 => x"08081c1c",
   972 => x"7c181000",
   973 => x"0010187c",
   974 => x"7c301000",
   975 => x"0010307c",
   976 => x"60603010",
   977 => x"00061e78",
   978 => x"183c6642",
   979 => x"0042663c",
   980 => x"c26a3878",
   981 => x"00386cc6",
   982 => x"60000060",
   983 => x"00600000",
   984 => x"5c5b5e0e",
   985 => x"86fc0e5d",
   986 => x"d1c17e71",
   987 => x"c04cbfd0",
   988 => x"c41ec04b",
   989 => x"c402ab66",
   990 => x"c24dc087",
   991 => x"754dc187",
   992 => x"ee49731e",
   993 => x"86c887e2",
   994 => x"ef49e0c0",
   995 => x"a4c487eb",
   996 => x"f0496a4a",
   997 => x"c9f187f2",
   998 => x"c184cc87",
   999 => x"abb7c883",
  1000 => x"87cdff04",
  1001 => x"4d268efc",
  1002 => x"4b264c26",
  1003 => x"711e4f26",
  1004 => x"d4d1c14a",
  1005 => x"d4d1c15a",
  1006 => x"4978c748",
  1007 => x"2687e1fe",
  1008 => x"1e731e4f",
  1009 => x"b7c04a71",
  1010 => x"87d303aa",
  1011 => x"bfdcccc1",
  1012 => x"c187c405",
  1013 => x"c087c24b",
  1014 => x"e0ccc14b",
  1015 => x"c187c45b",
  1016 => x"fc5ae0cc",
  1017 => x"dcccc148",
  1018 => x"c14a78bf",
  1019 => x"a2c0c19a",
  1020 => x"87e7ec49",
  1021 => x"4f264b26",
  1022 => x"c44a711e",
  1023 => x"49721e66",
  1024 => x"fc87f1eb",
  1025 => x"1e4f268e",
  1026 => x"c348d4ff",
  1027 => x"d0ff78ff",
  1028 => x"78e1c048",
  1029 => x"c148d4ff",
  1030 => x"c4487178",
  1031 => x"08d4ff30",
  1032 => x"48d0ff78",
  1033 => x"2678e0c0",
  1034 => x"5b5e0e4f",
  1035 => x"ec0e5d5c",
  1036 => x"48a6c886",
  1037 => x"c47e78c0",
  1038 => x"78bfec80",
  1039 => x"d1c180f8",
  1040 => x"e878bfd0",
  1041 => x"ccc14cbf",
  1042 => x"e349bfdc",
  1043 => x"eecb87fb",
  1044 => x"87cccb49",
  1045 => x"c758a6d4",
  1046 => x"87efe749",
  1047 => x"c9059870",
  1048 => x"4966cc87",
  1049 => x"c10299c1",
  1050 => x"66d087c4",
  1051 => x"ec7ec14d",
  1052 => x"ccc14bbf",
  1053 => x"e349bfdc",
  1054 => x"497587cf",
  1055 => x"7087edca",
  1056 => x"87d70298",
  1057 => x"bfc4ccc1",
  1058 => x"c1b9c149",
  1059 => x"7159c8cc",
  1060 => x"cb87f4fd",
  1061 => x"c7ca49ee",
  1062 => x"c74d7087",
  1063 => x"87ebe649",
  1064 => x"ff059870",
  1065 => x"497387c7",
  1066 => x"fe0599c1",
  1067 => x"026e87ff",
  1068 => x"c187e3c0",
  1069 => x"4abfdccc",
  1070 => x"ccc1bac1",
  1071 => x"0afc5ae0",
  1072 => x"9ac10a7a",
  1073 => x"49a2c0c1",
  1074 => x"c187d0e9",
  1075 => x"fae549da",
  1076 => x"48a6c887",
  1077 => x"ccc178c1",
  1078 => x"c105bfdc",
  1079 => x"c0c887c5",
  1080 => x"ccc14dc0",
  1081 => x"49134bc8",
  1082 => x"87dfe549",
  1083 => x"c2029870",
  1084 => x"c1b47587",
  1085 => x"ff052db7",
  1086 => x"497487ec",
  1087 => x"7199ffc3",
  1088 => x"fb49c01e",
  1089 => x"497487f2",
  1090 => x"7129b7c8",
  1091 => x"fb49c11e",
  1092 => x"86c887e6",
  1093 => x"e449fdc3",
  1094 => x"fac387f1",
  1095 => x"87ebe449",
  1096 => x"7487d4c7",
  1097 => x"99ffc349",
  1098 => x"712cb7c8",
  1099 => x"029c74b4",
  1100 => x"ccc187df",
  1101 => x"c749bfd8",
  1102 => x"987087f2",
  1103 => x"87c4c005",
  1104 => x"87d34cc0",
  1105 => x"c749e0c2",
  1106 => x"ccc187d6",
  1107 => x"c6c058dc",
  1108 => x"d8ccc187",
  1109 => x"7478c048",
  1110 => x"0599c849",
  1111 => x"c387cec0",
  1112 => x"e6e349f5",
  1113 => x"c2497087",
  1114 => x"e7c00299",
  1115 => x"d4d1c187",
  1116 => x"cac002bf",
  1117 => x"88c14887",
  1118 => x"58d8d1c1",
  1119 => x"c487d0c0",
  1120 => x"e0c14a66",
  1121 => x"c0026a82",
  1122 => x"ff4b87c5",
  1123 => x"c80f7349",
  1124 => x"78c148a6",
  1125 => x"99c44974",
  1126 => x"87cec005",
  1127 => x"e249f2c3",
  1128 => x"497087e9",
  1129 => x"c00299c2",
  1130 => x"d1c187f0",
  1131 => x"487ebfd4",
  1132 => x"03a8b7c7",
  1133 => x"6e87cbc0",
  1134 => x"c180c148",
  1135 => x"c058d8d1",
  1136 => x"66c487d3",
  1137 => x"80e0c148",
  1138 => x"bf6e7e70",
  1139 => x"87c5c002",
  1140 => x"7349fe4b",
  1141 => x"48a6c80f",
  1142 => x"fdc378c1",
  1143 => x"87ebe149",
  1144 => x"99c24970",
  1145 => x"87e9c002",
  1146 => x"bfd4d1c1",
  1147 => x"87c9c002",
  1148 => x"48d4d1c1",
  1149 => x"d3c078c0",
  1150 => x"4866c487",
  1151 => x"7080e0c1",
  1152 => x"02bf6e7e",
  1153 => x"4b87c5c0",
  1154 => x"0f7349fd",
  1155 => x"c148a6c8",
  1156 => x"49fac378",
  1157 => x"7087f4e0",
  1158 => x"0299c249",
  1159 => x"c187edc0",
  1160 => x"48bfd4d1",
  1161 => x"03a8b7c7",
  1162 => x"c187c9c0",
  1163 => x"c748d4d1",
  1164 => x"87d3c078",
  1165 => x"c14866c4",
  1166 => x"7e7080e0",
  1167 => x"c002bf6e",
  1168 => x"fc4b87c5",
  1169 => x"c80f7349",
  1170 => x"78c148a6",
  1171 => x"d1c17ec0",
  1172 => x"50c048cc",
  1173 => x"c349eecb",
  1174 => x"a6d487c6",
  1175 => x"ccd1c158",
  1176 => x"c105bf97",
  1177 => x"497487de",
  1178 => x"0599f0c3",
  1179 => x"c187cdc0",
  1180 => x"dfff49da",
  1181 => x"987087d5",
  1182 => x"87c8c102",
  1183 => x"bfe87ec1",
  1184 => x"ffc3494b",
  1185 => x"2bb7c899",
  1186 => x"ccc1b371",
  1187 => x"ff49bfdc",
  1188 => x"d087f6da",
  1189 => x"d3c24966",
  1190 => x"02987087",
  1191 => x"c187c6c0",
  1192 => x"c148ccd1",
  1193 => x"ccd1c150",
  1194 => x"c005bf97",
  1195 => x"497387d6",
  1196 => x"0599f0c3",
  1197 => x"c187c5ff",
  1198 => x"deff49da",
  1199 => x"987087cd",
  1200 => x"87f8fe05",
  1201 => x"e0c0026e",
  1202 => x"48a6cc87",
  1203 => x"bfd4d1c1",
  1204 => x"4966cc78",
  1205 => x"66c491cc",
  1206 => x"70807148",
  1207 => x"02bf6e7e",
  1208 => x"4b87c6c0",
  1209 => x"734966cc",
  1210 => x"0266c80f",
  1211 => x"c187c8c0",
  1212 => x"49bfd4d1",
  1213 => x"ec87e9f1",
  1214 => x"264d268e",
  1215 => x"264b264c",
  1216 => x"0000004f",
  1217 => x"00000000",
  1218 => x"14111258",
  1219 => x"231c1b1d",
  1220 => x"9491595a",
  1221 => x"f4ebf2f5",
  1222 => x"00000000",
  1223 => x"00000000",
  1224 => x"ff4a711e",
  1225 => x"7249bfc8",
  1226 => x"4f2648a1",
  1227 => x"bfc8ff1e",
  1228 => x"c0c0fe89",
  1229 => x"a9c0c0c0",
  1230 => x"c087c401",
  1231 => x"c187c24a",
  1232 => x"2648724a",
  1233 => x"00085f4f",
  1234 => x"00085f00",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
